//-----------------------------------------------------------------------------------
// CRC module for data[127:0] , crc[15:0]=1+x^5+x^12+x^16, reset active low 0x0000
//-----------------------------------------------------------------------------------
module crc_cacul(
  input [127:0] data_to_crc,
  input crc16_valid,
  output [15:0] data_from_crc,
  input rst_n,
  input clk_in
  output crc16_ready
  );

  reg [15:0] lfsr_q,lfsr_c;
  reg crc16_ready;

  assign data_from_crc = lfsr_q;

  always @(*) begin
    lfsr_c[0] = lfsr_q[1] ^ lfsr_q[3] ^ lfsr_q[6] ^ lfsr_q[9] ^ lfsr_q[11] ^ lfsr_q[15] ^ data_to_crc[0] ^ data_to_crc[4] ^ data_to_crc[8] ^ data_to_crc[11] ^ data_to_crc[12] ^ data_to_crc[19] ^ data_to_crc[20] ^ data_to_crc[22] ^ data_to_crc[26] ^ data_to_crc[27] ^ data_to_crc[28] ^ data_to_crc[32] ^ data_to_crc[33] ^ data_to_crc[35] ^ data_to_crc[42] ^ data_to_crc[48] ^ data_to_crc[49] ^ data_to_crc[51] ^ data_to_crc[52] ^ data_to_crc[55] ^ data_to_crc[56] ^ data_to_crc[58] ^ data_to_crc[63] ^ data_to_crc[64] ^ data_to_crc[65] ^ data_to_crc[66] ^ data_to_crc[67] ^ data_to_crc[70] ^ data_to_crc[72] ^ data_to_crc[74] ^ data_to_crc[75] ^ data_to_crc[77] ^ data_to_crc[80] ^ data_to_crc[81] ^ data_to_crc[82] ^ data_to_crc[84] ^ data_to_crc[86] ^ data_to_crc[88] ^ data_to_crc[95] ^ data_to_crc[96] ^ data_to_crc[98] ^ data_to_crc[104] ^ data_to_crc[106] ^ data_to_crc[107] ^ data_to_crc[108] ^ data_to_crc[109] ^ data_to_crc[110] ^ data_to_crc[113] ^ data_to_crc[115] ^ data_to_crc[118] ^ data_to_crc[121] ^ data_to_crc[123] ^ data_to_crc[127];
    lfsr_c[1] = lfsr_q[2] ^ lfsr_q[4] ^ lfsr_q[7] ^ lfsr_q[10] ^ lfsr_q[12] ^ data_to_crc[1] ^ data_to_crc[5] ^ data_to_crc[9] ^ data_to_crc[12] ^ data_to_crc[13] ^ data_to_crc[20] ^ data_to_crc[21] ^ data_to_crc[23] ^ data_to_crc[27] ^ data_to_crc[28] ^ data_to_crc[29] ^ data_to_crc[33] ^ data_to_crc[34] ^ data_to_crc[36] ^ data_to_crc[43] ^ data_to_crc[49] ^ data_to_crc[50] ^ data_to_crc[52] ^ data_to_crc[53] ^ data_to_crc[56] ^ data_to_crc[57] ^ data_to_crc[59] ^ data_to_crc[64] ^ data_to_crc[65] ^ data_to_crc[66] ^ data_to_crc[67] ^ data_to_crc[68] ^ data_to_crc[71] ^ data_to_crc[73] ^ data_to_crc[75] ^ data_to_crc[76] ^ data_to_crc[78] ^ data_to_crc[81] ^ data_to_crc[82] ^ data_to_crc[83] ^ data_to_crc[85] ^ data_to_crc[87] ^ data_to_crc[89] ^ data_to_crc[96] ^ data_to_crc[97] ^ data_to_crc[99] ^ data_to_crc[105] ^ data_to_crc[107] ^ data_to_crc[108] ^ data_to_crc[109] ^ data_to_crc[110] ^ data_to_crc[111] ^ data_to_crc[114] ^ data_to_crc[116] ^ data_to_crc[119] ^ data_to_crc[122] ^ data_to_crc[124];
    lfsr_c[2] = lfsr_q[0] ^ lfsr_q[3] ^ lfsr_q[5] ^ lfsr_q[8] ^ lfsr_q[11] ^ lfsr_q[13] ^ data_to_crc[2] ^ data_to_crc[6] ^ data_to_crc[10] ^ data_to_crc[13] ^ data_to_crc[14] ^ data_to_crc[21] ^ data_to_crc[22] ^ data_to_crc[24] ^ data_to_crc[28] ^ data_to_crc[29] ^ data_to_crc[30] ^ data_to_crc[34] ^ data_to_crc[35] ^ data_to_crc[37] ^ data_to_crc[44] ^ data_to_crc[50] ^ data_to_crc[51] ^ data_to_crc[53] ^ data_to_crc[54] ^ data_to_crc[57] ^ data_to_crc[58] ^ data_to_crc[60] ^ data_to_crc[65] ^ data_to_crc[66] ^ data_to_crc[67] ^ data_to_crc[68] ^ data_to_crc[69] ^ data_to_crc[72] ^ data_to_crc[74] ^ data_to_crc[76] ^ data_to_crc[77] ^ data_to_crc[79] ^ data_to_crc[82] ^ data_to_crc[83] ^ data_to_crc[84] ^ data_to_crc[86] ^ data_to_crc[88] ^ data_to_crc[90] ^ data_to_crc[97] ^ data_to_crc[98] ^ data_to_crc[100] ^ data_to_crc[106] ^ data_to_crc[108] ^ data_to_crc[109] ^ data_to_crc[110] ^ data_to_crc[111] ^ data_to_crc[112] ^ data_to_crc[115] ^ data_to_crc[117] ^ data_to_crc[120] ^ data_to_crc[123] ^ data_to_crc[125];
    lfsr_c[3] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[4] ^ lfsr_q[6] ^ lfsr_q[9] ^ lfsr_q[12] ^ lfsr_q[14] ^ data_to_crc[3] ^ data_to_crc[7] ^ data_to_crc[11] ^ data_to_crc[14] ^ data_to_crc[15] ^ data_to_crc[22] ^ data_to_crc[23] ^ data_to_crc[25] ^ data_to_crc[29] ^ data_to_crc[30] ^ data_to_crc[31] ^ data_to_crc[35] ^ data_to_crc[36] ^ data_to_crc[38] ^ data_to_crc[45] ^ data_to_crc[51] ^ data_to_crc[52] ^ data_to_crc[54] ^ data_to_crc[55] ^ data_to_crc[58] ^ data_to_crc[59] ^ data_to_crc[61] ^ data_to_crc[66] ^ data_to_crc[67] ^ data_to_crc[68] ^ data_to_crc[69] ^ data_to_crc[70] ^ data_to_crc[73] ^ data_to_crc[75] ^ data_to_crc[77] ^ data_to_crc[78] ^ data_to_crc[80] ^ data_to_crc[83] ^ data_to_crc[84] ^ data_to_crc[85] ^ data_to_crc[87] ^ data_to_crc[89] ^ data_to_crc[91] ^ data_to_crc[98] ^ data_to_crc[99] ^ data_to_crc[101] ^ data_to_crc[107] ^ data_to_crc[109] ^ data_to_crc[110] ^ data_to_crc[111] ^ data_to_crc[112] ^ data_to_crc[113] ^ data_to_crc[116] ^ data_to_crc[118] ^ data_to_crc[121] ^ data_to_crc[124] ^ data_to_crc[126];
    lfsr_c[4] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[2] ^ lfsr_q[5] ^ lfsr_q[7] ^ lfsr_q[10] ^ lfsr_q[13] ^ lfsr_q[15] ^ data_to_crc[4] ^ data_to_crc[8] ^ data_to_crc[12] ^ data_to_crc[15] ^ data_to_crc[16] ^ data_to_crc[23] ^ data_to_crc[24] ^ data_to_crc[26] ^ data_to_crc[30] ^ data_to_crc[31] ^ data_to_crc[32] ^ data_to_crc[36] ^ data_to_crc[37] ^ data_to_crc[39] ^ data_to_crc[46] ^ data_to_crc[52] ^ data_to_crc[53] ^ data_to_crc[55] ^ data_to_crc[56] ^ data_to_crc[59] ^ data_to_crc[60] ^ data_to_crc[62] ^ data_to_crc[67] ^ data_to_crc[68] ^ data_to_crc[69] ^ data_to_crc[70] ^ data_to_crc[71] ^ data_to_crc[74] ^ data_to_crc[76] ^ data_to_crc[78] ^ data_to_crc[79] ^ data_to_crc[81] ^ data_to_crc[84] ^ data_to_crc[85] ^ data_to_crc[86] ^ data_to_crc[88] ^ data_to_crc[90] ^ data_to_crc[92] ^ data_to_crc[99] ^ data_to_crc[100] ^ data_to_crc[102] ^ data_to_crc[108] ^ data_to_crc[110] ^ data_to_crc[111] ^ data_to_crc[112] ^ data_to_crc[113] ^ data_to_crc[114] ^ data_to_crc[117] ^ data_to_crc[119] ^ data_to_crc[122] ^ data_to_crc[125] ^ data_to_crc[127];
    lfsr_c[5] = lfsr_q[0] ^ lfsr_q[2] ^ lfsr_q[8] ^ lfsr_q[9] ^ lfsr_q[14] ^ lfsr_q[15] ^ data_to_crc[0] ^ data_to_crc[4] ^ data_to_crc[5] ^ data_to_crc[8] ^ data_to_crc[9] ^ data_to_crc[11] ^ data_to_crc[12] ^ data_to_crc[13] ^ data_to_crc[16] ^ data_to_crc[17] ^ data_to_crc[19] ^ data_to_crc[20] ^ data_to_crc[22] ^ data_to_crc[24] ^ data_to_crc[25] ^ data_to_crc[26] ^ data_to_crc[28] ^ data_to_crc[31] ^ data_to_crc[35] ^ data_to_crc[37] ^ data_to_crc[38] ^ data_to_crc[40] ^ data_to_crc[42] ^ data_to_crc[47] ^ data_to_crc[48] ^ data_to_crc[49] ^ data_to_crc[51] ^ data_to_crc[52] ^ data_to_crc[53] ^ data_to_crc[54] ^ data_to_crc[55] ^ data_to_crc[57] ^ data_to_crc[58] ^ data_to_crc[60] ^ data_to_crc[61] ^ data_to_crc[64] ^ data_to_crc[65] ^ data_to_crc[66] ^ data_to_crc[67] ^ data_to_crc[68] ^ data_to_crc[69] ^ data_to_crc[71] ^ data_to_crc[74] ^ data_to_crc[79] ^ data_to_crc[81] ^ data_to_crc[84] ^ data_to_crc[85] ^ data_to_crc[87] ^ data_to_crc[88] ^ data_to_crc[89] ^ data_to_crc[91] ^ data_to_crc[93] ^ data_to_crc[95] ^ data_to_crc[96] ^ data_to_crc[98] ^ data_to_crc[100] ^ data_to_crc[101] ^ data_to_crc[103] ^ data_to_crc[104] ^ data_to_crc[106] ^ data_to_crc[107] ^ data_to_crc[108] ^ data_to_crc[110] ^ data_to_crc[111] ^ data_to_crc[112] ^ data_to_crc[114] ^ data_to_crc[120] ^ data_to_crc[121] ^ data_to_crc[126] ^ data_to_crc[127];
    lfsr_c[6] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[3] ^ lfsr_q[9] ^ lfsr_q[10] ^ lfsr_q[15] ^ data_to_crc[1] ^ data_to_crc[5] ^ data_to_crc[6] ^ data_to_crc[9] ^ data_to_crc[10] ^ data_to_crc[12] ^ data_to_crc[13] ^ data_to_crc[14] ^ data_to_crc[17] ^ data_to_crc[18] ^ data_to_crc[20] ^ data_to_crc[21] ^ data_to_crc[23] ^ data_to_crc[25] ^ data_to_crc[26] ^ data_to_crc[27] ^ data_to_crc[29] ^ data_to_crc[32] ^ data_to_crc[36] ^ data_to_crc[38] ^ data_to_crc[39] ^ data_to_crc[41] ^ data_to_crc[43] ^ data_to_crc[48] ^ data_to_crc[49] ^ data_to_crc[50] ^ data_to_crc[52] ^ data_to_crc[53] ^ data_to_crc[54] ^ data_to_crc[55] ^ data_to_crc[56] ^ data_to_crc[58] ^ data_to_crc[59] ^ data_to_crc[61] ^ data_to_crc[62] ^ data_to_crc[65] ^ data_to_crc[66] ^ data_to_crc[67] ^ data_to_crc[68] ^ data_to_crc[69] ^ data_to_crc[70] ^ data_to_crc[72] ^ data_to_crc[75] ^ data_to_crc[80] ^ data_to_crc[82] ^ data_to_crc[85] ^ data_to_crc[86] ^ data_to_crc[88] ^ data_to_crc[89] ^ data_to_crc[90] ^ data_to_crc[92] ^ data_to_crc[94] ^ data_to_crc[96] ^ data_to_crc[97] ^ data_to_crc[99] ^ data_to_crc[101] ^ data_to_crc[102] ^ data_to_crc[104] ^ data_to_crc[105] ^ data_to_crc[107] ^ data_to_crc[108] ^ data_to_crc[109] ^ data_to_crc[111] ^ data_to_crc[112] ^ data_to_crc[113] ^ data_to_crc[115] ^ data_to_crc[121] ^ data_to_crc[122] ^ data_to_crc[127];
    lfsr_c[7] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[2] ^ lfsr_q[4] ^ lfsr_q[10] ^ lfsr_q[11] ^ data_to_crc[2] ^ data_to_crc[6] ^ data_to_crc[7] ^ data_to_crc[10] ^ data_to_crc[11] ^ data_to_crc[13] ^ data_to_crc[14] ^ data_to_crc[15] ^ data_to_crc[18] ^ data_to_crc[19] ^ data_to_crc[21] ^ data_to_crc[22] ^ data_to_crc[24] ^ data_to_crc[26] ^ data_to_crc[27] ^ data_to_crc[28] ^ data_to_crc[30] ^ data_to_crc[33] ^ data_to_crc[37] ^ data_to_crc[39] ^ data_to_crc[40] ^ data_to_crc[42] ^ data_to_crc[44] ^ data_to_crc[49] ^ data_to_crc[50] ^ data_to_crc[51] ^ data_to_crc[53] ^ data_to_crc[54] ^ data_to_crc[55] ^ data_to_crc[56] ^ data_to_crc[57] ^ data_to_crc[59] ^ data_to_crc[60] ^ data_to_crc[62] ^ data_to_crc[63] ^ data_to_crc[66] ^ data_to_crc[67] ^ data_to_crc[68] ^ data_to_crc[69] ^ data_to_crc[70] ^ data_to_crc[71] ^ data_to_crc[73] ^ data_to_crc[76] ^ data_to_crc[81] ^ data_to_crc[83] ^ data_to_crc[86] ^ data_to_crc[87] ^ data_to_crc[89] ^ data_to_crc[90] ^ data_to_crc[91] ^ data_to_crc[93] ^ data_to_crc[95] ^ data_to_crc[97] ^ data_to_crc[98] ^ data_to_crc[100] ^ data_to_crc[102] ^ data_to_crc[103] ^ data_to_crc[105] ^ data_to_crc[106] ^ data_to_crc[108] ^ data_to_crc[109] ^ data_to_crc[110] ^ data_to_crc[112] ^ data_to_crc[113] ^ data_to_crc[114] ^ data_to_crc[116] ^ data_to_crc[122] ^ data_to_crc[123];
    lfsr_c[8] = lfsr_q[1] ^ lfsr_q[2] ^ lfsr_q[3] ^ lfsr_q[5] ^ lfsr_q[11] ^ lfsr_q[12] ^ data_to_crc[3] ^ data_to_crc[7] ^ data_to_crc[8] ^ data_to_crc[11] ^ data_to_crc[12] ^ data_to_crc[14] ^ data_to_crc[15] ^ data_to_crc[16] ^ data_to_crc[19] ^ data_to_crc[20] ^ data_to_crc[22] ^ data_to_crc[23] ^ data_to_crc[25] ^ data_to_crc[27] ^ data_to_crc[28] ^ data_to_crc[29] ^ data_to_crc[31] ^ data_to_crc[34] ^ data_to_crc[38] ^ data_to_crc[40] ^ data_to_crc[41] ^ data_to_crc[43] ^ data_to_crc[45] ^ data_to_crc[50] ^ data_to_crc[51] ^ data_to_crc[52] ^ data_to_crc[54] ^ data_to_crc[55] ^ data_to_crc[56] ^ data_to_crc[57] ^ data_to_crc[58] ^ data_to_crc[60] ^ data_to_crc[61] ^ data_to_crc[63] ^ data_to_crc[64] ^ data_to_crc[67] ^ data_to_crc[68] ^ data_to_crc[69] ^ data_to_crc[70] ^ data_to_crc[71] ^ data_to_crc[72] ^ data_to_crc[74] ^ data_to_crc[77] ^ data_to_crc[82] ^ data_to_crc[84] ^ data_to_crc[87] ^ data_to_crc[88] ^ data_to_crc[90] ^ data_to_crc[91] ^ data_to_crc[92] ^ data_to_crc[94] ^ data_to_crc[96] ^ data_to_crc[98] ^ data_to_crc[99] ^ data_to_crc[101] ^ data_to_crc[103] ^ data_to_crc[104] ^ data_to_crc[106] ^ data_to_crc[107] ^ data_to_crc[109] ^ data_to_crc[110] ^ data_to_crc[111] ^ data_to_crc[113] ^ data_to_crc[114] ^ data_to_crc[115] ^ data_to_crc[117] ^ data_to_crc[123] ^ data_to_crc[124];
    lfsr_c[9] = lfsr_q[0] ^ lfsr_q[2] ^ lfsr_q[3] ^ lfsr_q[4] ^ lfsr_q[6] ^ lfsr_q[12] ^ lfsr_q[13] ^ data_to_crc[4] ^ data_to_crc[8] ^ data_to_crc[9] ^ data_to_crc[12] ^ data_to_crc[13] ^ data_to_crc[15] ^ data_to_crc[16] ^ data_to_crc[17] ^ data_to_crc[20] ^ data_to_crc[21] ^ data_to_crc[23] ^ data_to_crc[24] ^ data_to_crc[26] ^ data_to_crc[28] ^ data_to_crc[29] ^ data_to_crc[30] ^ data_to_crc[32] ^ data_to_crc[35] ^ data_to_crc[39] ^ data_to_crc[41] ^ data_to_crc[42] ^ data_to_crc[44] ^ data_to_crc[46] ^ data_to_crc[51] ^ data_to_crc[52] ^ data_to_crc[53] ^ data_to_crc[55] ^ data_to_crc[56] ^ data_to_crc[57] ^ data_to_crc[58] ^ data_to_crc[59] ^ data_to_crc[61] ^ data_to_crc[62] ^ data_to_crc[64] ^ data_to_crc[65] ^ data_to_crc[68] ^ data_to_crc[69] ^ data_to_crc[70] ^ data_to_crc[71] ^ data_to_crc[72] ^ data_to_crc[73] ^ data_to_crc[75] ^ data_to_crc[78] ^ data_to_crc[83] ^ data_to_crc[85] ^ data_to_crc[88] ^ data_to_crc[89] ^ data_to_crc[91] ^ data_to_crc[92] ^ data_to_crc[93] ^ data_to_crc[95] ^ data_to_crc[97] ^ data_to_crc[99] ^ data_to_crc[100] ^ data_to_crc[102] ^ data_to_crc[104] ^ data_to_crc[105] ^ data_to_crc[107] ^ data_to_crc[108] ^ data_to_crc[110] ^ data_to_crc[111] ^ data_to_crc[112] ^ data_to_crc[114] ^ data_to_crc[115] ^ data_to_crc[116] ^ data_to_crc[118] ^ data_to_crc[124] ^ data_to_crc[125];
    lfsr_c[10] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[3] ^ lfsr_q[4] ^ lfsr_q[5] ^ lfsr_q[7] ^ lfsr_q[13] ^ lfsr_q[14] ^ data_to_crc[5] ^ data_to_crc[9] ^ data_to_crc[10] ^ data_to_crc[13] ^ data_to_crc[14] ^ data_to_crc[16] ^ data_to_crc[17] ^ data_to_crc[18] ^ data_to_crc[21] ^ data_to_crc[22] ^ data_to_crc[24] ^ data_to_crc[25] ^ data_to_crc[27] ^ data_to_crc[29] ^ data_to_crc[30] ^ data_to_crc[31] ^ data_to_crc[33] ^ data_to_crc[36] ^ data_to_crc[40] ^ data_to_crc[42] ^ data_to_crc[43] ^ data_to_crc[45] ^ data_to_crc[47] ^ data_to_crc[52] ^ data_to_crc[53] ^ data_to_crc[54] ^ data_to_crc[56] ^ data_to_crc[57] ^ data_to_crc[58] ^ data_to_crc[59] ^ data_to_crc[60] ^ data_to_crc[62] ^ data_to_crc[63] ^ data_to_crc[65] ^ data_to_crc[66] ^ data_to_crc[69] ^ data_to_crc[70] ^ data_to_crc[71] ^ data_to_crc[72] ^ data_to_crc[73] ^ data_to_crc[74] ^ data_to_crc[76] ^ data_to_crc[79] ^ data_to_crc[84] ^ data_to_crc[86] ^ data_to_crc[89] ^ data_to_crc[90] ^ data_to_crc[92] ^ data_to_crc[93] ^ data_to_crc[94] ^ data_to_crc[96] ^ data_to_crc[98] ^ data_to_crc[100] ^ data_to_crc[101] ^ data_to_crc[103] ^ data_to_crc[105] ^ data_to_crc[106] ^ data_to_crc[108] ^ data_to_crc[109] ^ data_to_crc[111] ^ data_to_crc[112] ^ data_to_crc[113] ^ data_to_crc[115] ^ data_to_crc[116] ^ data_to_crc[117] ^ data_to_crc[119] ^ data_to_crc[125] ^ data_to_crc[126];
    lfsr_c[11] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[2] ^ lfsr_q[4] ^ lfsr_q[5] ^ lfsr_q[6] ^ lfsr_q[8] ^ lfsr_q[14] ^ lfsr_q[15] ^ data_to_crc[6] ^ data_to_crc[10] ^ data_to_crc[11] ^ data_to_crc[14] ^ data_to_crc[15] ^ data_to_crc[17] ^ data_to_crc[18] ^ data_to_crc[19] ^ data_to_crc[22] ^ data_to_crc[23] ^ data_to_crc[25] ^ data_to_crc[26] ^ data_to_crc[28] ^ data_to_crc[30] ^ data_to_crc[31] ^ data_to_crc[32] ^ data_to_crc[34] ^ data_to_crc[37] ^ data_to_crc[41] ^ data_to_crc[43] ^ data_to_crc[44] ^ data_to_crc[46] ^ data_to_crc[48] ^ data_to_crc[53] ^ data_to_crc[54] ^ data_to_crc[55] ^ data_to_crc[57] ^ data_to_crc[58] ^ data_to_crc[59] ^ data_to_crc[60] ^ data_to_crc[61] ^ data_to_crc[63] ^ data_to_crc[64] ^ data_to_crc[66] ^ data_to_crc[67] ^ data_to_crc[70] ^ data_to_crc[71] ^ data_to_crc[72] ^ data_to_crc[73] ^ data_to_crc[74] ^ data_to_crc[75] ^ data_to_crc[77] ^ data_to_crc[80] ^ data_to_crc[85] ^ data_to_crc[87] ^ data_to_crc[90] ^ data_to_crc[91] ^ data_to_crc[93] ^ data_to_crc[94] ^ data_to_crc[95] ^ data_to_crc[97] ^ data_to_crc[99] ^ data_to_crc[101] ^ data_to_crc[102] ^ data_to_crc[104] ^ data_to_crc[106] ^ data_to_crc[107] ^ data_to_crc[109] ^ data_to_crc[110] ^ data_to_crc[112] ^ data_to_crc[113] ^ data_to_crc[114] ^ data_to_crc[116] ^ data_to_crc[117] ^ data_to_crc[118] ^ data_to_crc[120] ^ data_to_crc[126] ^ data_to_crc[127];
    lfsr_c[12] = lfsr_q[2] ^ lfsr_q[5] ^ lfsr_q[7] ^ lfsr_q[11] ^ data_to_crc[0] ^ data_to_crc[4] ^ data_to_crc[7] ^ data_to_crc[8] ^ data_to_crc[15] ^ data_to_crc[16] ^ data_to_crc[18] ^ data_to_crc[22] ^ data_to_crc[23] ^ data_to_crc[24] ^ data_to_crc[28] ^ data_to_crc[29] ^ data_to_crc[31] ^ data_to_crc[38] ^ data_to_crc[44] ^ data_to_crc[45] ^ data_to_crc[47] ^ data_to_crc[48] ^ data_to_crc[51] ^ data_to_crc[52] ^ data_to_crc[54] ^ data_to_crc[59] ^ data_to_crc[60] ^ data_to_crc[61] ^ data_to_crc[62] ^ data_to_crc[63] ^ data_to_crc[66] ^ data_to_crc[68] ^ data_to_crc[70] ^ data_to_crc[71] ^ data_to_crc[73] ^ data_to_crc[76] ^ data_to_crc[77] ^ data_to_crc[78] ^ data_to_crc[80] ^ data_to_crc[82] ^ data_to_crc[84] ^ data_to_crc[91] ^ data_to_crc[92] ^ data_to_crc[94] ^ data_to_crc[100] ^ data_to_crc[102] ^ data_to_crc[103] ^ data_to_crc[104] ^ data_to_crc[105] ^ data_to_crc[106] ^ data_to_crc[109] ^ data_to_crc[111] ^ data_to_crc[114] ^ data_to_crc[117] ^ data_to_crc[119] ^ data_to_crc[123];
    lfsr_c[13] = lfsr_q[0] ^ lfsr_q[3] ^ lfsr_q[6] ^ lfsr_q[8] ^ lfsr_q[12] ^ data_to_crc[1] ^ data_to_crc[5] ^ data_to_crc[8] ^ data_to_crc[9] ^ data_to_crc[16] ^ data_to_crc[17] ^ data_to_crc[19] ^ data_to_crc[23] ^ data_to_crc[24] ^ data_to_crc[25] ^ data_to_crc[29] ^ data_to_crc[30] ^ data_to_crc[32] ^ data_to_crc[39] ^ data_to_crc[45] ^ data_to_crc[46] ^ data_to_crc[48] ^ data_to_crc[49] ^ data_to_crc[52] ^ data_to_crc[53] ^ data_to_crc[55] ^ data_to_crc[60] ^ data_to_crc[61] ^ data_to_crc[62] ^ data_to_crc[63] ^ data_to_crc[64] ^ data_to_crc[67] ^ data_to_crc[69] ^ data_to_crc[71] ^ data_to_crc[72] ^ data_to_crc[74] ^ data_to_crc[77] ^ data_to_crc[78] ^ data_to_crc[79] ^ data_to_crc[81] ^ data_to_crc[83] ^ data_to_crc[85] ^ data_to_crc[92] ^ data_to_crc[93] ^ data_to_crc[95] ^ data_to_crc[101] ^ data_to_crc[103] ^ data_to_crc[104] ^ data_to_crc[105] ^ data_to_crc[106] ^ data_to_crc[107] ^ data_to_crc[110] ^ data_to_crc[112] ^ data_to_crc[115] ^ data_to_crc[118] ^ data_to_crc[120] ^ data_to_crc[124];
    lfsr_c[14] = lfsr_q[1] ^ lfsr_q[4] ^ lfsr_q[7] ^ lfsr_q[9] ^ lfsr_q[13] ^ data_to_crc[2] ^ data_to_crc[6] ^ data_to_crc[9] ^ data_to_crc[10] ^ data_to_crc[17] ^ data_to_crc[18] ^ data_to_crc[20] ^ data_to_crc[24] ^ data_to_crc[25] ^ data_to_crc[26] ^ data_to_crc[30] ^ data_to_crc[31] ^ data_to_crc[33] ^ data_to_crc[40] ^ data_to_crc[46] ^ data_to_crc[47] ^ data_to_crc[49] ^ data_to_crc[50] ^ data_to_crc[53] ^ data_to_crc[54] ^ data_to_crc[56] ^ data_to_crc[61] ^ data_to_crc[62] ^ data_to_crc[63] ^ data_to_crc[64] ^ data_to_crc[65] ^ data_to_crc[68] ^ data_to_crc[70] ^ data_to_crc[72] ^ data_to_crc[73] ^ data_to_crc[75] ^ data_to_crc[78] ^ data_to_crc[79] ^ data_to_crc[80] ^ data_to_crc[82] ^ data_to_crc[84] ^ data_to_crc[86] ^ data_to_crc[93] ^ data_to_crc[94] ^ data_to_crc[96] ^ data_to_crc[102] ^ data_to_crc[104] ^ data_to_crc[105] ^ data_to_crc[106] ^ data_to_crc[107] ^ data_to_crc[108] ^ data_to_crc[111] ^ data_to_crc[113] ^ data_to_crc[116] ^ data_to_crc[119] ^ data_to_crc[121] ^ data_to_crc[125];
    lfsr_c[15] = lfsr_q[0] ^ lfsr_q[2] ^ lfsr_q[5] ^ lfsr_q[8] ^ lfsr_q[10] ^ lfsr_q[14] ^ data_to_crc[3] ^ data_to_crc[7] ^ data_to_crc[10] ^ data_to_crc[11] ^ data_to_crc[18] ^ data_to_crc[19] ^ data_to_crc[21] ^ data_to_crc[25] ^ data_to_crc[26] ^ data_to_crc[27] ^ data_to_crc[31] ^ data_to_crc[32] ^ data_to_crc[34] ^ data_to_crc[41] ^ data_to_crc[47] ^ data_to_crc[48] ^ data_to_crc[50] ^ data_to_crc[51] ^ data_to_crc[54] ^ data_to_crc[55] ^ data_to_crc[57] ^ data_to_crc[62] ^ data_to_crc[63] ^ data_to_crc[64] ^ data_to_crc[65] ^ data_to_crc[66] ^ data_to_crc[69] ^ data_to_crc[71] ^ data_to_crc[73] ^ data_to_crc[74] ^ data_to_crc[76] ^ data_to_crc[79] ^ data_to_crc[80] ^ data_to_crc[81] ^ data_to_crc[83] ^ data_to_crc[85] ^ data_to_crc[87] ^ data_to_crc[94] ^ data_to_crc[95] ^ data_to_crc[97] ^ data_to_crc[103] ^ data_to_crc[105] ^ data_to_crc[106] ^ data_to_crc[107] ^ data_to_crc[108] ^ data_to_crc[109] ^ data_to_crc[112] ^ data_to_crc[114] ^ data_to_crc[117] ^ data_to_crc[120] ^ data_to_crc[122] ^ data_to_crc[126];

  end // always

  always @(posedge clk_in or negedge rst_n) begin
    if(!rst_n) begin
      lfsr_q <= {16{1'b0}};
    end
    else begin
        if(crc16_valid) begin
          lfsr_q <= lfsr_c;
          crc16_ready <= 1'b1;
        end
        else begin
          lfsr_q <= lfsr_q;
          crc16_ready <= 1'b0;
        end
    end
  end // always
endmodule // crc